/****************************************************************************
 * Convert.sv
 ****************************************************************************/

/**
 * Module: Convert
 * 
 * TODO: Add module documentation
 */
module Convert(		maxnum,
					SCnum,
					clk,
					Bnum);
	
	
	


endmodule


