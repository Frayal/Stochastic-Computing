/****************************************************************************
 * Clock.sv
 ****************************************************************************/

/**
 * Module: Clock
 * 
 * TODO: Add module documentation
 */
module Clock;


endmodule


