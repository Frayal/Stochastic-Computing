/****************************************************************************
 * addition.sv
 ****************************************************************************/

/**
 * Module: addition
 * 
 * TODO: Add module documentation
 */
module addition;


endmodule


