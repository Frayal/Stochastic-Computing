/****************************************************************************
 * Convert.sv
 ****************************************************************************/

/**
 * Module: Convert
 * 
 * TODO: Add module documentation
 */
module Convert;


endmodule


